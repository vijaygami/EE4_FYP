** Profile: "SCHEMATIC1-fitting"  [ C:\Users\Vijay\Google Drive\PSpice\FYP\Intro\Fitting\fitting-pspicefiles\schematic1\fitting.sim ] 

** Creating circuit file "fitting.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../fitting-pspicefiles/vteam.lib" 
* From [PSPICE NETLIST] section of C:\Users\Vijay\Documents\PSpice\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 7.95s 0 0.05m SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
