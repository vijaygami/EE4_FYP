** Profile: "SCHEMATIC1-imply_gate"  [ C:\Users\Vijay\Google Drive\PSpice\FYP\MAGIC\NOR\imply_gate-pspicefiles\schematic1\imply_gate.sim ] 

** Creating circuit file "imply_gate.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../imply_gate-pspicefiles/vteam.lib" 
.LIB "../../../imply_gate-pspicefiles/imply_gate.lib" 
* From [PSPICE NETLIST] section of C:\Users\Vijay\Documents\PSpice\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 320 0 30m SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
