** Profile: "SCHEMATIC1-Initial_investigations"  [ C:\Users\Vijay\Google Drive\PSpice\FYP\Intro\heuristic_threshold\initial_investigations-pspicefiles\schematic1\initial_investigations.sim ] 

** Creating circuit file "Initial_investigations.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../initial_investigations-pspicefiles/vteam.lib" 
.LIB "../../../initial_investigations-pspicefiles/team.lib" 
* From [PSPICE NETLIST] section of C:\Users\Vijay\Documents\PSpice\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1010 1000 2m SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
