** Profile: "SCHEMATIC1-bias"  [ C:\Users\Vijay\Google Drive\PSpice\FYP\MRL\xor_buf\gates-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../gates-pspicefiles/gates.lib" 
.LIB "../../../gates-pspicefiles/vteam.lib" 
* From [PSPICE NETLIST] section of C:\Users\Vijay\Documents\PSpice\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 79.99 0 10m SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
