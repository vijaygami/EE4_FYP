** Profile: "SCHEMATIC1-xor_unbuf"  [ C:\Users\Vijay\Google Drive\PSpice\FYP\MRL\xor_unbuf\xor_unbuf-pspicefiles\schematic1\xor_unbuf.sim ] 

** Creating circuit file "xor_unbuf.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../xor_unbuf-pspicefiles/vteam.lib" 
.LIB "../../../xor_unbuf-pspicefiles/xor_unbuf.lib" 
* From [PSPICE NETLIST] section of C:\Users\Vijay\Documents\PSpice\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 79.99 0 10m SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
