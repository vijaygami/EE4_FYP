** Profile: "SCHEMATIC1-memrist_intro"  [ C:\Users\Vijay\Google Drive\PSpice\FYP\Intro\memrist_intro\memrst_intro-pspicefiles\schematic1\memrist_intro.sim ] 

** Creating circuit file "memrist_intro.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../memrst_intro-pspicefiles/team.lib" 
.LIB "../../../memrst_intro-pspicefiles/vteam.lib" 
* From [PSPICE NETLIST] section of C:\Users\Vijay\Documents\PSpice\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1s 0 0.005m SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
